`define channel_num 4
//hls�㷨Ԥ�� decode��������Ӧ�ô�ԼΪdecode���ʵ�2/3-3/4
//��Ҫ�ǿ�InvMixColumns((state_t*)in);